`timescale 1ns / 1ns

module Depacketizer (
    
);

    

endmodule
